** sch_path: /home/tare/Desktop/Analog design/dff.sch
**.subckt dff
V4 D GND pulse(0 VDD {TCLK/4} TRF TRF {3*TCLK} {4*TCLK})
.save i(v4)
V5 CLK GND pulse(0 VDD 0 TRF TRF {TCLK/2} TCLK)
.save i(v5)
V3 RST GND pulse(0 VDD {3.5*TCLK} TRF TRF {2*TCLK} {16*TCLK})
.save i(v3)
V1 SET GND pulse(0 VDD {11.5*TCLK} TRF TRF {2*TCLK} {16*TCLK})
.save i(v1)
C1 Q GND 1P m=1
C2 QB GND 1P m=1
**** begin user architecture code



*These are the values of the parameters to be used
.param VDD=2 VCC=VDD
.param TRF=1n TCLK=100n
.param TSTOP={20*TCLK} TDROP=0
*Analysis setup and control statements
.tran 100p {TSTOP} {TDROP}
*save all voltages and currents
.save all
*options for an accurate precision output
.options reltol=1e-6 vntol=1u abstol=1p
* option to make output file ascii
*.options filetype=ascii




a3 D CLK SET RST Q QB my_dff
.model my_dff d_dff(clk_delay = 0.5e-9 set_delay = 0.5e-9                    rreset_delay = 0.5e-9
+ ic = 0 rise_delay = 0.5e-9  fall_delay = 0.5e-9)


**** end user architecture code
**.ends
.GLOBAL GND
.end
