** sch_path: /home/tare/Desktop/Analog design/inv_tb.sch
**.subckt inv_tb
V1 A GND pulse(0 VDD 0 TRF TRF {TCLK/2} TCLK)
.save i(v1)
C1 Y GND 100f m=1
**** begin user architecture code



*These are the values of the parameters to be used
.param VDD=2 VCC=VDD
.param TRF=1n TCLK=100n
.param TSTOP={5*TCLK} TDROP=0
*Analysis setup and control statements
.tran 100p {TSTOP} {TDROP}
*save all voltages and currents
.save all
*options for an accurate precision output
.options reltol=1e-6 vntol=1u abstol=1p
* option to make output file ascii
*.options filetype=ascii




a1 A Y inv1
.model inv1 d_inverter(rise_delay = 0.5e-9 fall_delay = 0.5e-9  input_load = 0.1e-12)


**** end user architecture code
**.ends
.GLOBAL GND
.end
